library verilog;
use verilog.vl_types.all;
entity testbench_SHIFT_LEFT is
end testbench_SHIFT_LEFT;
