library verilog;
use verilog.vl_types.all;
entity testbench_ALU_3 is
end testbench_ALU_3;
