library verilog;
use verilog.vl_types.all;
entity testbench_SHIFT_LEFT_LOGIC is
end testbench_SHIFT_LEFT_LOGIC;
