library verilog;
use verilog.vl_types.all;
entity testebench_ADDER_FULL is
end testebench_ADDER_FULL;
